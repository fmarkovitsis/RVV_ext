module tb;
  reg 
